module adder(input [31:0] inp1 , inp2,output reg [31:0] out);
	assign out = inp1 + inp2;
endmodule
